../../../dmem/hdl/sv/dmem.sv