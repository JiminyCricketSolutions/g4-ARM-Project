../../../alu/hdl/sv/alu.sv