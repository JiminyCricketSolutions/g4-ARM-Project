../../../datapath/hdl/sv/datapath.sv