../../../adder/hdl/sv/adder.sv