../../../condlogic/hdl/sv/condlogic.sv