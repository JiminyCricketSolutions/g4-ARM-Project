../../../ram/hdl/sv/ram.sv