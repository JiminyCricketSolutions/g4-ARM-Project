../../../main_decoder/hdl/sv/decoder.sv