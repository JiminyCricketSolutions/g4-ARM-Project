../../../extend/hdl/sv/extender.sv