../../../controller/hdl/sv/controller.sv