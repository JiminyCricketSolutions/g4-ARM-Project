../../../mux2/hdl/sv/mux2.sv