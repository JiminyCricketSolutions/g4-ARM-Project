../../../flopenr/hdl/sv/flopenr.sv