../../../condcheck/hdl/sv/condcheck.sv