../../../imem/hdl/sv/imem.sv