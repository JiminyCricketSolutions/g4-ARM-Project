../../../ARM-single-cycle/hdl/sv/ARMSC.sv