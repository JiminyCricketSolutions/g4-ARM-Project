../../../registerfile/hdl/sv/registerfile.sv