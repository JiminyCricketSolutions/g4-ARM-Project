../../../flopr/hdl/sv/flopr.sv